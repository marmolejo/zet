`timescale 1ns/10ps

module ram_2k_attr (clk, rst, cs, we, addr, rdata, wdata);
  // IO Ports
  input clk;
  input rst;
  input cs;
  input we;
  input [10:0] addr;
  output [7:0] rdata;
  input [7:0] wdata;

  // Net declarations
  wire dp;
  wire rw;

  // Module instantiations
  RAMB16_S9 ram (.DO(rdata),
                 .DOP (dp),
                 .ADDR (addr),
                 .CLK (clk),
                 .DI (wdata),
                 .DIP (dp),
                 .EN (cs),
                 .SSR (rst),
                 .WE (rw));

    defparam ram.INIT_00 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_01 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_02 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_03 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_04 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_05 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_06 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_07 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_08 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_09 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_0A = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_0B = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_0C = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_0D = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_0E = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_0F = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_10 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_11 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_12 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_13 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_14 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_15 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_16 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_17 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_18 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_19 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_1A = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_1B = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_1C = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_1D = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_1E = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_1F = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_20 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_21 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_22 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_23 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_24 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_25 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_26 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_27 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_28 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_29 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_2A = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_2B = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_2C = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_2D = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_2E = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_2F = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_30 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_31 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_32 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_33 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_34 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_35 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_36 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_37 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_38 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_39 = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_3A = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_3B = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_3C = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_3D = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_3E = 256'h0707070707070707070707070707070707070707070707070707070707070707;
    defparam ram.INIT_3F = 256'h0707070707070707070707070707070707070707070707070707070707070707;

  // Assignments
  assign rw = ~we;
endmodule